Journal||(?:[\t ]*@HEADER_DOC_JOURNAL)[\t ]+
Title||(?:[\t ]*@HEADER_DOC_TITLE)[\t ]+
Abstract||(?:[\t ]*@HEADER_DOC_ABSTRACT)[\t ]+
Summary||(?:[\t ]*@HEADER_DOC_SUMMARY)[\t ]+
Inclusion Criteria||(?:[\t ]*@HEADER_DOC_INCLUSION_CRITERIA)[\t ]+
Exclusion Criteria||(?:[\t ]*@HEADER_DOC_EXCLUSION_CRITERIA)[\t ]+
Unknown Criteria||(?:[\t ]*@HEADER_DOC_UNKNOWN_CRITERIA)[\t ]+
Mesh Terms||(?:[\t ]*@HEADER_DOC_MESH_TERMS)[\t ]+
Primary Outcomes||(?:[\t ]*@HEADER_DOC_PRIMARY_OUTCOMES)[\t ]+
Secondary Outcomes||(?:[\t ]*@HEADER_DOC_SECONDARY_OUTCOMES)[\t ]+
